//
// SPDX-FileCopyrightText: Copyright 2023-2024 Darryl Miles
// SPDX-License-Identifier: Apache2.0
//

//
//

// One of these is expected to be set by the synthesis environment:
// `define TECH_SKY130 1
// `define TECH_IHP130 1
// `define TECH_FPGA 1

// Defined when running project in Vivado/Xilinx/Arty-A7
//`define FPGA_XILINX_7SERIES 1
